library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity toplevel_tb is
end entity;

architecture toplevel_tb_arch of toplevel_tb is
    
end architecture;